p, q, p^q, !q&p, !(p&q)